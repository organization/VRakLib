module vraklib

struct Packet {
    buffer byteptr
}