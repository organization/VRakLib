module raklib

struct RakLib {
    server_ip string
    server_port u16

    running bool
}