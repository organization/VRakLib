module vraklib

struct Packet {

}