module vraklib

struct VRakLib {
    server_ip string
    server_port u16

    running bool
}