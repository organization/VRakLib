module raklib

struct Packet {

}