module vraklib

struct LoginPaket {
    packet Packet
}